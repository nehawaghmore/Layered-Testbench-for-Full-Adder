class transaction;

// Stimulus are declared with rand keyword
 
  rand bit in1;  
  rand bit in2;
  rand bit cin;
  
  bit sum;
  bit cout; 
endclass
